module  tft_pic
(
    input   wire            tft_clk     ,
    input   wire            sys_rst_n   ,
    input   wire    [9:0]   pix_x       ,
    input   wire    [9:0]   pix_y       ,
    
    output  reg     [15:0]  pix_data       

);

parameter   CHAR_B_H = 112,
            CHAR_B_V = 104;
            
parameter   CHAR_W = 256,
            CHAR_H = 64;
            
parameter   BLACK  = 16'h0000,
            GOLDEN = 16'hFEC0;

wire    [9:0]   char_x  ;
wire    [9:0]   char_y  ;
reg     [255:0] char    [63:0];
//二位寄存器数组，描述存储器结构
//定义一个存储器，地址为0~63，每个存储单元都是256比特
//与一维的reg变量不同的是，不可对存储单元进行位选择或部分选择
//可以为每个存储单元单独赋值
//一维： reg [3:0] char;  位选择 char[1] = 1; 部分选择 char[1:0] = 2'b10

assign  char_x = (((pix_x >= CHAR_B_H) && (pix_x < CHAR_B_H + CHAR_W)) &&
                  ((pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H))) 
                  ? (pix_x - CHAR_B_H) : 10'h3ff;

assign  char_y = (((pix_x >= CHAR_B_H) && (pix_x < CHAR_B_H + CHAR_W)) &&
                 ((pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H)))  
                  ? (pix_y - CHAR_B_V) : 10'h3ff;
       
always@(posedge tft_clk)                  
    begin
        char[ 0]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[ 1]    <=  256'h00001E0000000000000000000000000000000000000000000000000000000000;
        char[ 2]    <=  256'h000002000003F000000000000000000000000000000000000000000000000000;
        char[ 3]    <=  256'h0003E30026020800000000000000000000000000000000000000000000000000;
        char[ 4]    <=  256'h0000E3003383E830060000000000000000000000000000000000000000000000;
        char[ 5]    <=  256'h0000630010826818C20000000000000000000000000000000000000000000000;
        char[ 6]    <=  256'h071C633010824808410000000000000000000000000000000000000000000000;
        char[ 7]    <=  256'h019463C010831808210000000000000000000000000000000000000000000000;
        char[ 8]    <=  256'h019C6300117FF8082F0000000000000000000000000000000000000000000000;
        char[ 9]    <=  256'h0100FFC013860818610000000000000000000000000000000000000000000000;  
        char[10]    <=  256'h07F8FFFC10041033FF0000000000000000000000000000000000000000000000;
        char[11]    <=  256'h00004000000030FC010000000000000000000400000000000000000000000000;
        char[12]    <=  256'h0000000000003000000000000000000000000600000000000080000000000000;
        char[13]    <=  256'h000000000000100000000000000000000000037F700000000080000000100000;
        char[14]    <=  256'h0000000000000000000000000000000000000180478000000080000000100000;
        char[15]    <=  256'h00000007FFFFF000017E00000000000000000080408000000080000000100000;
        char[16]    <=  256'h00000002000000000100A0000000000000000083C18000000000000386100000;
        char[17]    <=  256'h00000001C000000001000800000000C100000043C3000000008000023F100000;
        char[18]    <=  256'h007FF001C000000001000100000000C100000027C601F8000200000101100000;
        char[19]    <=  256'h01C01E01C0000000000000C0000001230000003FDC0010000480000001800000;
        char[20]    <=  256'h07000300C000000001000020006F822200000010B00060000000000100D00000;
        char[21]    <=  256'h0C000101C0000000000000100280020400000000000080000000000001000000;
        char[22]    <=  256'h18003901C0000000010000080C00041800000000800100000480000001920000;
        char[23]    <=  256'h13800102C000000000000008200000180000000080060000080040008F820000;
        char[24]    <=  256'h2000790140000000010000184000100000000000000C00000001800070110000;
        char[25]    <=  256'h27C0F101C0000000000000308000202400000000000700000803000035550000;
        char[26]    <=  256'h6780F103800000000000002100000002000000008000C00109080000401C0000;
        char[27]    <=  256'h400001038000000001000043000000800000000000002001C020000000300000;
        char[28]    <=  256'h40000301800000000000008200008002000000010000F3603080000041D00000;
        char[29]    <=  256'h4008020780000000000003040000000100000000007F88181600000007000000;  
        char[30]    <=  256'h401802038000000000000804000002008000000100600F8819000000A8000000;
        char[31]    <=  256'h40380207F00000000100100800011ED4FF700000004008E80700003D20200000;
        char[32]    <=  256'h40380203EFDA000000008008001EBFFFFFF00007004008380700000080000000;
        char[33]    <=  256'h40080207000FF000000900080004004A4940000DC040080006000002E0000000;
        char[34]    <=  256'h400006030000000000A000100003EA00400DE009602000000200000820400000;
        char[35]    <=  256'h4000440700000001DA000010000000004000000820200800020001A030000000;
        char[36]    <=  256'h2000C40200000000000000100209000020000009600008000900030030400000;
        char[37]    <=  256'h2181840600000000000000100200000020000009C01000000100060008000000;
        char[38]    <=  256'h30F70C0600000000000000100202000030000005001008000080000034400000;
        char[39]    <=  256'h101C080600000000020000100620000010000007000800000080000046000000;  
        char[40]    <=  256'h1800100600000000000000000A08000010000009000008001000000003C00000;
        char[41]    <=  256'h0C00200400000000000000100A40000010000025000408000040000121800000;
        char[42]    <=  256'h0601C00600000000020000101250000010000085000000000020000000800000;
        char[43]    <=  256'h03FF0006000000000000001022A0000018000203000210004000000420800000;
        char[44]    <=  256'h000000060000000000000010C2C0000018002803000010002010000000800000;
        char[45]    <=  256'h0000000E0000000002000011028000000002C003000110000010002020800000;
        char[46]    <=  256'h0000000E000000000000000E0280000000070002000010010008000042800000;
        char[47]    <=  256'h0000000E0000000000000000020000000000A442000091C00000000062C60000;
        char[48]    <=  256'h0000000C000000000400000000000000000000044220D9324004020065060000;
        char[49]    <=  256'h0000000C00000000000000000000000000000000000050000004000069060000;  
        char[50]    <=  256'h0000000C0000000000000000000000000000000000003004800408002FC60000;
        char[51]    <=  256'h00000008000000000400000000000000000000000000200000020000010E0000;
        char[52]    <=  256'h00000008000000000000000000000000000000000000000880036000013A0000;
        char[53]    <=  256'h0000000000000000000000000000000000000000000000110001C00000020000;
        char[54]    <=  256'h0000000000000000040000000000000000000000000000160000000001020000;
        char[55]    <=  256'h00000000000000000000000000000000000000000000001C0000000001170000;
        char[56]    <=  256'h000000000000000000000000000000000000000000000018000000000F770000;
        char[57]    <=  256'h0000000000000000040000000000000000000000000000000000000033820000;
        char[58]    <=  256'h000000000000000000000000000000000000000000000000000000001F7C0000;
        char[59]    <=  256'h000000000000000000000000000000000000000000000000000000000FF00000;  
        char[60]    <=  256'h0000000000000000040000000000000000000000000000000000000007060000;
        char[61]    <=  256'h0000000000000000040000000000000000000000000000000000000000030000;
        char[62]    <=  256'h0000000000000000040000000000000000000000000000000000000000000000;
        char[63]    <=  256'h0000000000000000040000000000000000000000000000000000000000000000;
  
    end 
                  
always@(posedge tft_clk or negedge sys_rst_n)                
    if(sys_rst_n == 1'b0)
        pix_data <= BLACK;
    else    if(((pix_x >= CHAR_B_H - 1'b1) && (pix_x < CHAR_B_H + CHAR_W - 1'b1)) &&  //提前一个时钟周期而不是提前一行
               ((pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H)) &&
               (char[char_y][10'd255 - char_x] == 1'b1))//防止左右颠倒
        pix_data <= GOLDEN;
    else
        pix_data <= BLACK;
                  
                  

endmodule