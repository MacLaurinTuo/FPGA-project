module  clk_gen(
    input   wire    inclk0  ,
    input   wire    arest   ,
    
    output  reg     c0

);







endmodule