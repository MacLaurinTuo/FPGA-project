module  vga_pic
(
    input   wire            vga_clk     ,
    input   wire            sys_rst_n   ,
    input   wire    [9:0]   pix_x       ,
    input   wire    [9:0]   pix_y       ,
    
    output  reg     [15:0]  pix_data       

);

parameter   CHAR_B_H = 192,
            CHAR_B_V = 208;
            
parameter   CHAR_W = 256,
            CHAR_H = 64;
            
parameter   BLACK  = 16'h0000,
            GOLDEN = 16'hFEC0;

wire    [9:0]   char_x  ;
wire    [9:0]   char_y  ;
reg     [255:0] char    [63:0];
//二位寄存器数组，描述存储器结构
//定义一个存储器，地址为0~63，每个存储单元都是256比特
//与一维的reg变量不同的是，不可对存储单元进行位选择或部分选择
//可以为每个存储单元单独赋值
//一维： reg [3:0] char;  位选择 char[1] = 1; 部分选择 char[1:0] = 2'b10

assign  char_x = (((pix_x >= CHAR_B_H) && (pix_x < CHAR_B_H + CHAR_W)) &&
                  ((pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H))) 
                  ? (pix_x - CHAR_B_H) : 10'h3ff;

assign  char_y = (((pix_x >= CHAR_B_H) && (pix_x < CHAR_B_H + CHAR_W)) &&
                 ((pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H)))  
                  ? (pix_y - CHAR_B_V) : 10'h3ff;
                  
always@(posedge vga_clk)                  
    begin
        char[ 0]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[ 1]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[ 2]    <=  256'h0000000000000000000000200000000000000000002000000008000010000000;
        char[ 3]    <=  256'h000000000000000000000038000000000000020000380000000600001C000000;
        char[ 4]    <=  256'h02000000000100000000003E0000000000000700003E0000000780001F000000;
        char[ 5]    <=  256'h03000070000380000000003E0000000000001F8000380000000700001E000000;
        char[ 6]    <=  256'h03FFFFF9FFFFE0000000003C000000000000FF8000380000000700001C000000;
        char[ 7]    <=  256'h0381C0708003E0000000003C00000000000FFC0000380000000700001C000000;
        char[ 8]    <=  256'h0381C070000780000000003C0000000000FFC00000380000000700001C000000;
        char[ 9]    <=  256'h0381C070000E00000000003C000000000F81C00000380000000700001C000000;   
        char[10]    <=  256'h0381C070001C00000000003C000000000001C00600380000000700001C000000;
        char[11]    <=  256'h0381C070303800000000003C000000000001C00380380000000700001C000000;
        char[12]    <=  256'h0381C070186000000000003C000000000001C001E0380000000700001C008000;
        char[13]    <=  256'h0381C0700E4000000000003C000000000001C000F038000000070C001C01C000;
        char[14]    <=  256'h0381C070078000000000003C000000000001C000F038000000071E801C03E000;
        char[15]    <=  256'h0381C07003C000000000003C001800000001C000783800001FFFFFFFFFFFF000;
        char[16]    <=  256'h03FFFFF001E000000000003C001C00000001C00030380000000700001C000000;
        char[17]    <=  256'h0381C07001F000000001003C003E00000001C00030380000000700001C000000;
        char[18]    <=  256'h0381C07000F000000003003C003F00000001C18000380000000700001C000000;
        char[19]    <=  256'h0381C070006040000002003C007C00000001C3C000380000000700001C000000;
        char[20]    <=  256'h0381C070006060000006003C00F800001FFFFFE000380000000700001C000000;
        char[21]    <=  256'h0381C0780000F0000006003C00F000000803C00000380000000700001C000000;
        char[22]    <=  256'h0381C077FFFFF8000006003C01E000000003C00000380000000700001C000000;
        char[23]    <=  256'h0381C07201C0F000000E003C03C000000003C00400380000000701001C060000;
        char[24]    <=  256'h0381C07001C1C000001E003C030000000007C00300380000000707801C0F0000;
        char[25]    <=  256'h0381C07001C18000003C003A060000000007C0038038000000073C7FFFFF8000;
        char[26]    <=  256'h03FFFFF001C30000007C007A0C000000000FE001E03800000007F008000F0000;
        char[27]    <=  256'h0381C07001C2000000F8007B18000000000FF800E0380000000FC00C000E0000;
        char[28]    <=  256'h0381C06001C6000001F8007930000000001FDE00F0380000003F0004001E0000;
        char[29]    <=  256'h0201C00001C0000001F00071E0000000001DCF007038000001FF0006001C0000;   
        char[30]    <=  256'h0001C00001C0000001E00071800000000039C780603860001FF70006001C0000;
        char[31]    <=  256'h0001C00001C00000000000F0C00000000039C3806038F0001FC7000200380000;
        char[32]    <=  256'h0001C00001C00000000000E0C00000000071C3800038F8000F07000300380000;
        char[33]    <=  256'h0001C02001C00000000000E0600000000061C180003FE0000407000300780000;
        char[34]    <=  256'h0001C07001C00000000001E07000000000E1C10000FC00000007000180700000;
        char[35]    <=  256'h0FFFC0F801C00000000001C03000000001C1C0003FB800000007000180E00000;
        char[36]    <=  256'h07FFFFFC01C00000000003C0380000000181C007F038000000070000C1E00000;
        char[37]    <=  256'h0001C00001C00000000003801C0000000301C0FE0038000000070000E1C00000;
        char[38]    <=  256'h0001C00001C00000000007800E0000000601C1C0003800000007000063C00000;
        char[39]    <=  256'h0001C00001C00000000007000F0000000C01C080003800000007000077800000;   
        char[40]    <=  256'h0001C00001C0000000000F00078000000801C00000380000000700003F000000;
        char[41]    <=  256'h0001C00001C0000000001E0003C000001001C00000380000000700003E000000;
        char[42]    <=  256'h0001C00001C0000000001C0003E000002001C00000380000000700003E000000;
        char[43]    <=  256'h0001C03E01C000000000380001F000000001C00000380000000700007F000000;
        char[44]    <=  256'h0001CFE001C000000000700000F800000001C0000038000000070000F7800000;
        char[45]    <=  256'h0003FE0001C000000000E000007E00000001C0000038000000070003E3E00000;
        char[46]    <=  256'h01FFE00001C000000003C000003F80000001C000003800000007000781F80000;
        char[47]    <=  256'h3FFE000001C0000000078000001FE0000001C000003800000E0F001F00FE0000;
        char[48]    <=  256'h1FE00001FFC00000000E0000000FFC000001C0000038000003FF007C003FE000;
        char[49]    <=  256'h1F0000003FC00000003C00000003F0000001C0000038000000FE01F0001FFC00;   
        char[50]    <=  256'h080000000F80000000F000000001C0000003C00000380000007E07800007E000;
        char[51]    <=  256'h000000000700000003C00000000080000003C00000380000001C1E000001C000;
        char[52]    <=  256'h00000000020000000E0000000000000000038000003800000010600000004000;
        char[53]    <=  256'h0000000000000000100000000000000000020000002000000000000000000000;
        char[54]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[55]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[56]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[57]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[58]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[59]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;   
        char[60]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[61]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[62]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[63]    <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
  
    end 
                  
always@(posedge vga_clk or negedge sys_rst_n)                
    if(sys_rst_n == 1'b0)
        pix_data <= BLACK;
    else    if(((pix_x >= CHAR_B_H - 1'b1) && (pix_x < CHAR_B_H + CHAR_W - 1'b1)) &&
               ((pix_y >= CHAR_B_V) && (pix_y < CHAR_B_V + CHAR_H)) &&
               (char[char_y][10'd256 - char_x] == 1'b1))//防止左右颠倒
        pix_data <= GOLDEN;
    else
        pix_data <= BLACK;
                  
                  

endmodule